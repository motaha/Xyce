Simple RC circuit
*.param Rval=1Meg Cval=100n sinfreq=1000 T1={Rval*Cval} Vval=12V T2={1/sinfreq}
.param Rval=1Meg Cval=100n sinfreq=1000 T1={Rval*Cval} Vval=1V T2={1/sinfreq}
Vsrc    1 0  DC 0V SIN(0V {Vval} {sinfreq} 0 0)
R1 1 2 {Rval}
C1 2 0 {Cval}
.print tran V(1) V(2) I(Vsrc)
.options timeint reltol=1e-4 abstol=1e-6 conststep=1 maxord=1
.options DEVICE voltlim=0
.tran 10us 300ms
.END
